`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 28.10.2025 11:50:44
// Design Name: 
// Module Name: testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1ns / 1ps

module testbench;
    reg [3:0] bcd_in;
    wire [3:0] excess3_out;

    BCD_2_EXCESS3 dut(bcd_in, excess3_out);

    always begin
        bcd_in= 4'd0;
    #10;
        bcd_in= 4'd1;
    #10;
        bcd_in= 4'd2;
    #10;
        bcd_in= 4'd3;
    #10;
        bcd_in= 4'd4;
    #10;
        bcd_in= 4'd5;
    #10;
        bcd_in= 4'd6;
    #10;
        bcd_in= 4'd7;
    #10;
        bcd_in= 4'd8;
    #10;
        bcd_in= 4'd9;
    #10;
        bcd_in= 4'd10;
    #10;
        bcd_in= 4'd11;
    #10;
        bcd_in= 4'd12;
    #10;
        bcd_in= 4'd13;
    #10;
        bcd_in= 4'd14;
    #10;
        bcd_in= 4'd15;
    #10;
    end
    
    initial begin
    $monitor("Input: %b  Excess-3 Code: %b", bcd_in, excess3_out);
    #160 $finish;
    end
endmodule
