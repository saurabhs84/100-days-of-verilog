`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08.12.2025 10:30:40
// Design Name: 
// Module Name: testbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module testbench;
parameter N=4;
reg clk,reset;
wire [N-1:0] gray;

Gray_Counter uut (.clk(clk),.reset(reset),.gray(gray));
always #5 clk=~clk;
initial begin
clk=0;
reset=1;#10
reset=0;
#100
reset=1;
#20
reset=0;
#200
$finish;
end
initial begin
$monitor("time=%t | clk=%b | reset=%b | gray=%b",$time,clk,reset,gray);
end
endmodule
